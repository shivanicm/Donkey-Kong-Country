module BananaAddr();

